module das68k();
endmodule
